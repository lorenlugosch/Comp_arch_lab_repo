-- Loren Lugosch
-- 260404057

-- Testbench for cache_SRAM.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY cache_SRAM_tb IS
END cache_SRAM_tb;

ARCHITECTURE behavior OF cache_SRAM_tb IS

...
END behavior;