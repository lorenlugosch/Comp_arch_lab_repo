-- Loren Lugosch
-- 260404057

-- This VHD describes a cache.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

-- cache entity adapted from given memory description entity --
ENTITY cache IS
	GENERIC(
		word_length : INTEGER := 32;
		address_length : INTEGER := 32;
		associativity : INTEGER := 1; --two-way associative?--
		index_length : INTEGER := 8; --256 cache lines means 8 bits of index--
		tag_length : INTEGER := 22; --32 address bits minus 10 = 22 tag bits--
		offset_length : INTEGER := 2; --4 words per line means 2 bits req'd to address a word--
		--SRAM_width : INTEGER := 150;
		number_of_cache_blocks : INTEGER := 256
	);
	PORT(
		clock : IN STD_LOGIC;
		writedata : IN STD_LOGIC_VECTOR (word_length-1 downto 0);
		addr : IN STD_LOGIC_VECTOR (31 downto 0);
		memwrite : IN STD_LOGIC;
		memread : IN STD_LOGIC;
		readdata : OUT STD_LOGIC_VECTOR (word_length-1 downto 0);
		waitrequest : OUT STD_LOGIC -- tells FSM to keep waiting--
	);
END cache;

ARCHITECTURE arch OF cache IS
  -- goes high when a read or write is requested by CPU --
  SIGNAL mem_request : STD_LOGIC;
  
	-- address decoding signals --
	SIGNAL input_tag : STD_LOGIC_VECTOR(tag_length-1 downto 0);
	SIGNAL input_index : INTEGER RANGE 0 to 255; --STD_LOGIC_VECTOR(index_length-1 downto 0); 
	SIGNAL input_offset : STD_LOGIC_VECTOR(1 downto 0);
	
	-- readdata for each word SRAM --
	SIGNAL readdata_zero : STD_LOGIC_VECTOR(word_length-1 downto 0);
	SIGNAL readdata_one : STD_LOGIC_VECTOR(word_length-1 downto 0);
	SIGNAL readdata_two : STD_LOGIC_VECTOR(word_length-1 downto 0);
	SIGNAL readdata_three : STD_LOGIC_VECTOR(word_length-1 downto 0);
	
	-- readdata for tag, dirty, valid --
	SIGNAL readdata_tag : STD_LOGIC_VECTOR(tag_length+2-1 downto 0);
	
	-- signals to make changes to tag/valid/dirty --
	SIGNAL writedata_tag : STD_LOGIC_VECTOR(tag_length+2-1 downto 0);
	
	-- signals for selecting a word to write to --
	SIGNAL memwrite_zero : STD_LOGIC;
	SIGNAL memwrite_one : STD_LOGIC;
	SIGNAL memwrite_two : STD_LOGIC;
	SIGNAL memwrite_three : STD_LOGIC;
	
	-- cache lines --
	COMPONENT cache_SRAM
		GENERIC (
			SRAM_width : INTEGER; -- \
			number_of_rows : INTEGER
		);
		PORT (
			clock : in STD_LOGIC;
			writedata : in STD_LOGIC_VECTOR(SRAM_width-1 downto 0);
			address : in INTEGER RANGE 0 to number_of_cache_blocks-1;
			writeenable : in STD_LOGIC;
			readdata : out STD_LOGIC_VECTOR(SRAM_width-1 downto 0)
		);
	END COMPONENT;
	
	BEGIN
	  -- detect memory access --
		mem_request <= memread or memwrite;
	  
	  -- decode address --
		input_tag <= addr(address_length-1 downto address_length-tag_length);
		input_index <= to_integer(unsigned(addr(address_length-tag_length-1 downto address_length-tag_length-index_length)));
		input_offset <= addr(offset_length-1 downto 0);
		
		-- select word to write --
		memwrite_zero <= memwrite and not input_offset(1) and not input_offset(0);
		memwrite_one <= memwrite and not input_offset(1) and input_offset(0);
		memwrite_two <= memwrite and input_offset(1) and not input_offset(0);
		memwrite_three <= memwrite and input_offset(1) and input_offset(0);
		
		-- tag SRAM contains: tag, dirty bit, valid bit
		tag_SRAM: cache_SRAM GENERIC MAP (SRAM_width => tag_length+2, number_of_rows => number_of_cache_blocks)
									PORT MAP (clock, writedata_tag, input_index, memwrite, readdata_tag);
		word_zero_SRAM: cache_SRAM GENERIC MAP (SRAM_width => word_length, number_of_rows => number_of_cache_blocks)
									PORT MAP (clock, writedata, input_index, memwrite_zero, readdata_zero);
		word_one_SRAM: cache_SRAM GENERIC MAP (SRAM_width => word_length, number_of_rows => number_of_cache_blocks)
									PORT MAP (clock, writedata, input_index, memwrite_one, readdata_one);
		word_two_SRAM: cache_SRAM GENERIC MAP (SRAM_width => word_length, number_of_rows => number_of_cache_blocks)
									PORT MAP (clock, writedata, input_index, memwrite_two, readdata_two);
		word_three_SRAM: cache_SRAM GENERIC MAP (SRAM_width => word_length, number_of_rows => number_of_cache_blocks)
									PORT MAP (clock, writedata, input_index, memwrite_three, readdata_three);
				
		-- "input_offset" represents which word of the cache line we want --
		-- use it to select which SRAM's output data we want to read --
		with input_offset select
			readdata <= readdata_zero when "00",
						   readdata_one when "01",
						   readdata_two when "10",
						   readdata_three when "11",
						   X"00000000" when others;
		
		-- dummy output to test address decoding --
		--readdata <= X"12345678";
		waitrequest <= '1';
	
END arch;