-- cache FSM