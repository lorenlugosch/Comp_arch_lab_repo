-- Loren Lugosch
-- 260404057
-- 
-- Out_FIFOs have a FIFO queue
-- connected to another router
-- in the network of cores
-- and an interface which tells 
-- the various in_FIFOs that 
-- they can write.
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.router_parameters.all;

entity out_FIFO is
	--generic ();
	--port ();
end out_FIFO;

architecture rtl of out_FIFO is

begin

end rtl;
